** sch_path: /home/juan/Documents/Workshop_ihp/Modulo_Analogico/Lab5/inverter/xschem/inverter.sch
.subckt inverter Vin VDD VSS Vout
*.PININFO Vin:I VDD:B VSS:B Vout:B
M1 Vout Vin VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=1
M2 Vout Vin VDD VDD sg13_lv_pmos w=3u l=1u ng=1 m=1
.ends
.end
