** sch_path: /home/juan/Documents/Workshop_ihp/Modulo_Analogico/Lab5/inverter/xschem/inverter_tb_tran.sch
**.subckt inverter_tb_tran
x1 Vin VDD VSS Vout inverter
C1 Vout VSS 100f m=1
V1 VSS GND 0
V2 VDD VSS 1.5
Vin Vin VSS PULSE(0 1.5 0 5n 5n 1u 2u)
**** begin user architecture code


.tran 1n 10u
.save all



.lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/juan/Documents/Workshop_ihp/Modulo_Analogico/Lab5/inverter/xschem/inverter.sym
** sch_path: /home/juan/Documents/Workshop_ihp/Modulo_Analogico/Lab5/inverter/xschem/inverter.sch
.subckt inverter Vin VDD VSS Vout
*.ipin Vin
*.iopin VDD
*.iopin VSS
*.iopin Vout
XM1 Vout Vin VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=1
XM2 Vout Vin VDD VDD sg13_lv_pmos w=3u l=1u ng=1 m=1
.ends

.GLOBAL GND
.end
